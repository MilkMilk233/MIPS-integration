`timescale 1ns/1ps

module alu_test;
reg[31:0] instruction,regA, regB;

wire[31:0] result;
wire[2:0] flags;

alu testalu(instruction,regA,regB, result, flags);

initial
begin

$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
$monitor("   %h:%h: %h :%h:%h:%h:  %b   :    %b     :    %b     :%b:%b:  %b",
instruction, testalu.opcode, testalu.func, regA ,regB, result, flags[2],flags[1],flags[0], testalu.rs_reg, testalu.rt_reg, testalu.reg_C);


//在本test sample里，rs对应regA（地址00000），rt对应regB（地址00001）


//add
// 3 + 9 = c
#10 instruction<=32'b000000_00000_00001_00011_00000_100000;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
$display("add");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
// 模拟溢出
#10 instruction<=32'b000000_00000_00001_00011_00000_100000;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
// 模拟溢出
#10 instruction<=32'b000000_00000_00001_00001_00000_100000;
regA<=32'b0100_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b0100_0000_0000_0000_0000_0000_0000_0001;
//相加等于0
#10 instruction<=32'b000000_00000_00001_00001_00000_100000;
regA<=32'b0000_0000_0000_0000_0000_0000_1101_1101;
regB<=32'b1111_1111_1111_1111_1111_1111_0010_0011;
//相加等于负数
#10 instruction<=32'b000000_00000_00001_00001_00000_100000;
regA<=32'b0000_0010_0010_0000_1000_1111_0101_1101;
regB<=32'b1111_1101_1101_1111_0111_0000_0010_0011;

//addi，这里是regA+imm sign extended
#10 instruction<=32'b001000_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_0000_0101_1100_0000_0001;
regB<=32'b1000_0000_0000_0101_1100_0101_1100_0001;
$display("addi");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001000_00000_00001_0000000000100010;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b1000_0000_0101_1100_0000_0000_0000_0001;

#10 instruction<=32'b001000_00000_00001_0000000000100000;
regA<=32'b1000_0000_0101_1100_0000_0000_0000_0001;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
//测试溢出
#10 instruction<=32'b001000_00000_00001_1111111111111111;
regA<=32'b0111_1111_1111_1111_0000_0000_0000_0001;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

//addu，本质上和add一样，由于不判断flags，故忽略
#10 instruction<=32'b000000_00000_00001_00001_00000_100001;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b0000_0000_0000_0101_1100_0000_0000_1001;
$display("addu");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_100001;
regA<=32'b1000_0000_0101_1100_0000_0000_0000_0001;
regB<=32'b1000_0000_0000_0101_1100_0000_0000_0001;

#10 instruction<=32'b000000_00000_00001_00001_00000_100001;
regA<=32'b0100_0000_0101_1100_0000_0000_0000_0001;
regB<=32'b0100_0000_0000_0101_1100_0000_0000_0001;

#10 instruction<=32'b000000_00000_00001_00001_00000_100001;
regA<=32'b0000_0000_0000_0000_0000_0000_1101_1101;
regB<=32'b1111_0101_1100_1111_1111_1111_0010_0011;

#10 instruction<=32'b000000_00000_00001_00001_00000_100001;
regA<=32'b0000_0000_0000_0101_1100_0000_0101_1101;
regB<=32'b1111_1111_0101_1100_1111_1111_0010_0011;

#10 instruction<=32'b000000_00000_00001_00001_00000_100001;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b0000_0101_1100_0000_0000_0000_0000_0000;

//addiu，本质上和addi一样，同上。
#10 instruction<=32'b001001_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
$display("addiu");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001001_00000_00001_1000000000100000;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b0000_0101_1100_0000_0000_0000_0000_0011;

#10 instruction<=32'b001001_00000_00001_0000000000000000;
regA<=32'b0000_0101_1100_0000_0000_0000_0000_0000;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//sub，用regA - regB
#10 instruction<=32'b000000_00000_00001_00001_00000_100010;
regA<=32'b1111_0000_0000_0000_0000_0000_0101_1101;
regB<=32'b0000_0101_1100_0000_0000_0000_0000_0001;
$display("sub");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_100010;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b0111_0000_0000_0000_0000_0000_0101_1101;

#10 instruction<=32'b000000_00000_00001_00001_00000_100010;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b1111_0000_0101_1100_0000_0101_1100_1101;

#10 instruction<=32'b000000_00000_00001_00001_00000_100010;
regA<=32'b0000_0000_0101_1100_0000_0000_0000_0000;
regB<=32'b0000_0000_0000_0000_0101_0101_1100_0000;

//subu，不考虑flags
#10 instruction<=32'b000000_00000_00001_00001_00000_100011;
regA<=32'b0111_0101_1100_0000_0101_1100_0101_1101;
regB<=32'b1000_0000_0000_1111_0000_0000_0000_0001;
$display("subu");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_100011;
regA<=32'b1000_0000_0000_1111_0000_0000_0000_0001;
regB<=32'b0111_0000_1111_0000_0000_0000_0101_1111;

#10 instruction<=32'b000000_00000_00001_00001_00000_100011;
regA<=32'b0000_0000_1111_0000_0000_0000_0000_0001;
regB<=32'b1111_0000_0000_0000_0000_0000_0101_0001;

#10 instruction<=32'b000000_00000_00001_00001_00000_100011;
regA<=32'b0000_0000_0000_0000_0000_1000_0000_1101;
regB<=32'b0000_0000_1111_0000_0000_0000_0101_1101;

#10 instruction<=32'b000000_00000_00001_00001_00000_100011;
regA<=32'b0000_0000_0000_0000_1111_0000_0000_0000;
regB<=32'b0000_1111_0000_1111_0000_0000_0000_0000;

//and
#10 instruction<=32'b000000_00000_00001_00001_00000_100100;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("and");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_100100;
regA<=32'b1000_0000_1001_0000_0000_0000_0000_0000;
regB<=32'b0000_0000_1001_0000_0000_0000_0011_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_100100;
regA<=32'b1000_1100_0010_0000_0000_0000_0000_0000;
regB<=32'b0100_0001_0000_0001_0110_0000_0011_1110;

#10 instruction<=32'b000000_00000_00001_00001_00000_100100;
regA<=32'b1000_0100_0100_1100_0000_0110_1100_0100;
regB<=32'b1111_1111_1100_0011_1101_1111_1111_1111;

//andi
#10 instruction<=32'b001100_00000_00001_1000000000100000;
regA<=32'b1000_0110_0000_0000_0000_0000_0000_0001;
regB<=32'b1000_0000_0110_0000_0000_0000_0000_0001;
$display("andi");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001100_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_0110_0000_0000_0010_0000;
regB<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 instruction<=32'b001100_00000_00001_1000000000100000;
regA<=32'b0000_0000_0000_0000_0110_0000_0000_0001;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//nor
#10 instruction<=32'b000000_00000_00001_00001_00000_100111;
regA<=32'b1000_0000_0010_0000_0000_0000_0000_0000;
regB<=32'b1111_1111_1101_1111_1111_1111_1111_1111;
$display("nor");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_100111;
regA<=32'b1000_0110_0000_0000_0000_0000_0000_0000;
regB<=32'b0000_0000_0000_1100_0000_0000_0011_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_100111;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

#10 instruction<=32'b000000_00000_00001_00001_00000_100111;
regA<=32'b1000_1100_1110_0000_1100_0000_0000_0000;
regB<=32'b0000_0010_0000_0000_0000_0000_0011_0010;

//or
#10 instruction<=32'b000000_00000_00001_00001_11000_100101;
regA<=32'b1111_1100_0010_1100_0010_0100_0100_0000;
regB<=32'b0000_0000_0000_1100_0100_0010_0001_0010;
$display("or");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_11000_100101;
regA<=32'b0100_0000_1111_1111_0000_0000_0010_0000;
regB<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

#10 instruction<=32'b000000_00000_00001_00001_11000_100101;
regA<=32'b0000_0000_0010_0100_0000_0000_0010_0000;
regB<=32'b0000_0000_1000_0100_0000_0000_0010_0000;

//ori
#10 instruction<=32'b001101_00000_00001_1000000000100000;
regA<=32'b1000_0000_1000_0010_0000_0000_0000_0001;
regB<=32'b1100_0000_0000_0010_0000_0000_0000_0001;
$display("ori");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001101_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_0100_0010_0001_0010_0000;
regB<=32'b1000_0000_0000_0100_0010_0001_1000_0001;

#10 instruction<=32'b001101_00000_00001_0000000000000000;
regA<=32'b0000_0000_0100_0000_0000_0000_0000_0000;
regB<=32'b0000_0000_1111_1111_0000_0000_0000_0011;

//xor
#10 instruction<=32'b000000_00000_00001_00001_00000_100110;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("xor");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_100110;
regA<=32'b1000_0000_0000_0010_0000_0000_0000_0000;
regB<=32'b0000_0000_1111_1111_0000_0000_0011_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_100110;
regA<=32'b1000_1100_0010_0010_0000_0010_0000_0000;
regB<=32'b0000_1111_1111_1000_0000_0000_0011_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_100110;
regA<=32'b1000_0000_0000_0000_0000_0010_0000_0000;
regB<=32'b1111_1111_1000_1011_1111_1111_1111_1111;

//xori
#10 instruction<=32'b001110_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_0000_0000_1000_1011_0001;
regB<=32'b1000_0000_1000_1011_0000_0000_1000_1011;
$display("xori");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001110_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_0100_0000_0000_0010_0000;
regB<=32'b1000_0000_0000_0100_0000_0010_0000_0001;

#10 instruction<=32'b001110_00000_00001_1000000000100000;
regA<=32'b0000_0000_0010_0000_0000_0111_0000_0001;
regB<=32'b0000_0000_1000_0000_0000_0010_0000_0011;

//beq/bne
#10 instruction<=32'b000101_00000_00001_1000000000100000;
regA<=32'b1000_0000_0100_0000_0000_0000_0000_0001;
regB<=32'b1000_0000_0100_0000_0000_0000_0000_0001;
$display("beq/bne");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000100_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_1000_0000_0000_0010_0000;
regB<=32'b1000_0000_0000_1000_0000_0000_0010_0000;

#10 instruction<=32'b000100_00000_00001_1000000000100000;
regA<=32'b0000_0000_0000_0010_0000_0000_0000_0001;
regB<=32'b0000_0000_0000_0010_0000_0000_0000_0001;

//slt
#10 instruction<=32'b000000_00000_00001_00001_00000_101010;
regA<=32'b1000_0000_0000_1000_1011_0000_0000_0000;
regB<=32'b1111_1000_1011_1111_1111_1111_1111_1111;
$display("slt");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_101010;
regA<=32'b1000_0000_1000_1011_0000_0000_0000_0000;
regB<=32'b0000_0000_0000_0000_0000_0000_0000_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_101010;
regA<=32'b0100_1100_0010_0000_0000_0000_0000_0000;
regB<=32'b0000_0000_0000_1000_1011_0000_0000_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_101010;
regA<=32'b1010_0000_0100_0000_0000_0000_0000_0000;
regB<=32'b1111_1111_1111_1011_1100_1000_1011_1111;

//slti
#10 instruction<=32'b001010_00000_00001_1000000000100000;
regA<=32'b1010_0000_0000_0000_0000_0000_0000_0001;
regB<=32'b1000_0000_0100_0000_0000_0000_1100_0001;
$display("slti");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001010_00000_00001_1000000000100000;
regA<=32'b1100_0000_1000_0000_0000_0000_0010_0000;
regB<=32'b1010_1000_0100_0000_0000_0110_0000_0001;

#10 instruction<=32'b001010_00000_00001_1000000000100000;
regA<=32'b0000_0000_1100_0100_0000_0000_0000_0001;
regB<=32'b0000_0110_0110_0010_0000_0110_0000_0011;

//sltu
#10 instruction<=32'b000000_00000_00001_00001_00000_101011;
regA<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
regB<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("sltu");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_00000_101011;
regA<=32'b1000_0000_0010_0000_0000_0000_1000_0000;
regB<=32'b0000_0000_0000_1111_1111_1111_1111_1111;

#10 instruction<=32'b000000_00000_00001_00001_00000_101011;
regA<=32'b1000_1100_0010_1100_0000_0000_0000_0000;
regB<=32'b0000_0110_1000_0000_0000_1100_0011_0010;

#10 instruction<=32'b000000_00000_00001_00001_00000_101011;
regA<=32'b1000_0000_1100_0000_0000_0000_0000_0000;
regB<=32'b1111_1111_1111_0011_1111_1111_1111_1111;

//stliu
#10 instruction<=32'b001011_00000_00001_0000000000100000;
regA<=32'b0000_0000_0000_0000_0100_0000_0000_0000;
regB<=32'b0000_0000_0000_0000_0000_0000_1000_0001;
$display("stliu");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b001011_00000_00001_0000000000010000;
regA<=32'b0000_0100_0000_0000_0100_0000_0010_0000;
regB<=32'b0000_0000_0100_0000_0000_0100_0000_0001;

#10 instruction<=32'b001011_00000_00001_1000000000100000;
regA<=32'b1000_0110_0000_0000_0000_0000_0000_0000;
regB<=32'b1000_0000_0000_0110_0000_0000_0000_1001;

#10 instruction<=32'b001011_00000_00001_1000000000100000;
regA<=32'b0100_0010_0000_0100_0000_0000_0000_0000;
regB<=32'b1000_0000_0100_0100_0110_0000_0000_0011;

//sw
#10 instruction<=32'b101011_00000_00001_1000000000100000;
regA<=32'b1100_0100_0000_0000_1100_0000_0000_0001;
regB<=32'b1010_0110_0000_0000_0000_1100_0000_0001;
$display("sw");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b101011_00000_00001_1000000000100000;
regA<=32'b1000_0000_0000_1100_0000_0000_0010_0000;
regB<=32'b1000_0000_0100_0000_0000_1111_0000_0001;

#10 instruction<=32'b101011_00000_00001_1000000000100000;
regA<=32'b0000_0000_0100_0000_1110_0000_0110_0001;
regB<=32'b0000_0110_0000_1100_0000_0000_0000_0011;

//lw
#10 instruction<=32'b100011_00000_00001_1000000000100000;
regA<=32'b1000_0000_0100_0000_0010_1100_0011_0001;
regB<=32'b1000_0110_0000_1100_0010_1100_1100_1101;
$display("lw");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b100011_00000_00001_1000000000100000;
regA<=32'b1000_0000_0010_0000_0010_0000_0010_0000;
regB<=32'b1000_0110_0000_0000_0000_0100_0000_0001;

#10 instruction<=32'b100011_00000_00001_1000000000100000;
regA<=32'b0000_0010_0010_0100_0000_0100_0000_0001;
regB<=32'b0000_0110_0000_1100_0000_0001_0000_0011;

//sll,将regB向左移动2位
#10 instruction<=32'b000000_00000_00001_00001_00010_000000;
regA<=32'b1111_1100_0010_0000_0000_0001_0000_0000;
regB<=32'b0000_0000_0000_0100_1010_0010_0000_0010;
$display("sll");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
//将regB向左移动24位
#10 instruction<=32'b000000_00000_00001_00001_11000_000000;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
regB<=32'b1111_0000_1111_0000_0000_1111_1111_1111;

//sllv,将regB向左移动regA位，填0
#10 instruction<=32'b000000_00000_00001_00001_11000_000100;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
regB<=32'b0000_0000_0000_0010_0100_0100_0010_0010;
$display("sllv");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_11000_000100;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
regB<=32'b0000_0000_1000_0101_0100_0000_0001_0000;

//srl，将regB向右移动2位，填0
#10 instruction<=32'b000000_00000_00001_00001_00010_000010;
regA<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
regB<=32'b1000_0010_0110_0110_1010_0110_0000_0010;
$display("srl");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_11000_000010;
regA<=32'b0100_0000_0000_0000_0000_0000_0000_0000;
regB<=32'b1111_0000_0000_0000_0000_0000_0000_0000;

//srlv，将regB向右移动2位，填0
#10 instruction<=32'b000000_00000_00001_00001_11000_000110;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
regB<=32'b1000_1010_0010_0100_1000_0100_0000_0010;
$display("srlv");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_11000_000110;
regA<=32'b1000_0000_0000_0000_0000_0000_0000_0010;
regB<=32'b0110_0010_0010_0000_0100_1101_0010_1000;

//sra，将regB向右移动2位，填msb
#10 instruction<=32'b000000_00000_00001_00001_00010_000011;
regA<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
regB<=32'b1000_0000_0000_0100_0010_0100_0100_0010;
$display("sra");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_11000_000011;
regA<=32'b0100_0000_0010_0000_0000_0000_0000_0000;
regB<=32'b1111_1001_1001_1111_0011_1111_0011_0000;

//srav，将regB向右移动2位,填msb
#10 instruction<=32'b000000_00000_00001_00001_11000_000111;
regA<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
regB<=32'b1000_0100_0100_1101_1100_0010_0010_0010;
$display("srav");
$display("instruction:op:func:  regA  :  regB  : result : zero : negative : overflow :               rs               :               rt               :            result_buffer");
#10 instruction<=32'b000000_00000_00001_00001_11000_000111;
regA<=32'b0000_0000_0100_0010_0001_0000_0000_0110;
regB<=32'b0100_0100_1100_1100_0000_0000_0101_0000;


#10 $finish;
end
endmodule